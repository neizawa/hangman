{"secret_word":"applicable","guessed_letters":["_","_","_","_","_","c","_","b","_","e"],"guess":11,"used_letters":["t","f","s","r","e","m","n","b","v","c","x"]}